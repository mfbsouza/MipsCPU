module Control (
	input clk,
);

endmodule: Control