module cpu(
	input clock,
	input reset,
	
);

logic meme [31:0]

Registrador Pc(
	//conexoes
);

Mux5 IorD(
	//conexoes
);

Memoria Mem(
	//conexoes
);

WriteMode WM(
	//conexoes
);

Registrador MDR(
	//conexoes
);

Instr_Reg IR(
	//conexoes
);

